`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    01:38:44 06/03/2021 
// Design Name: 
// Module Name:    RISC_TOP 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module RISC_TOP(input [31:0]A,B,input [15:0]ADD,input clk,rst,Asel, output [31:0]ALU_out,Data_out);


endmodule
